module cosrom (
	input c, // clock
	input [9:0] a0, a1, // angle
	output reg [34:0] d0, d1);

	reg [34:0] oreg0, oreg1;
	(* ram_style = "block" *) reg [34:0] bram[0:1023];

always @ (posedge c) begin
	oreg0 <= bram[a0];
	oreg1 <= bram[a1];
	d0 <= oreg0;
	d1 <= oreg1;
end

initial begin
	bram[0] <= 35'd34359730181;
	bram[1] <= 35'd34359689231;
	bram[2] <= 35'd34359566360;
	bram[3] <= 35'd34359369763;
	bram[4] <= 35'd34359083052;
	bram[5] <= 35'd34358722615;
	bram[6] <= 35'd34358272064;
	bram[7] <= 35'd34357747786;
	bram[8] <= 35'd34357141588;
	bram[9] <= 35'd34356453469;
	bram[10] <= 35'd34355691624;
	bram[11] <= 35'd34354839666;
	bram[12] <= 35'd34353905787;
	bram[13] <= 35'd34352898181;
	bram[14] <= 35'd34351808655;
	bram[15] <= 35'd34350637209;
	bram[16] <= 35'd34349383843;
	bram[17] <= 35'd34348048557;
	bram[18] <= 35'd34346631350;
	bram[19] <= 35'd34345140417;
	bram[20] <= 35'd34343559370;
	bram[21] <= 35'd34341904596;
	bram[22] <= 35'd34340167902;
	bram[23] <= 35'd34338349288;
	bram[24] <= 35'd34336448754;
	bram[25] <= 35'd34334466299;
	bram[26] <= 35'd34332410118;
	bram[27] <= 35'd34330263823;
	bram[28] <= 35'd34328043801;
	bram[29] <= 35'd34325741860;
	bram[30] <= 35'd34323349804;
	bram[31] <= 35'd34320892215;
	bram[32] <= 35'd34318344513;
	bram[33] <= 35'd34315714890;
	bram[34] <= 35'd34313011541;
	bram[35] <= 35'd34310218078;
	bram[36] <= 35'd34307350888;
	bram[37] <= 35'd34304401778;
	bram[38] <= 35'd34301370748;
	bram[39] <= 35'd34298257797;
	bram[40] <= 35'd34295071120;
	bram[41] <= 35'd34291794329;
	bram[42] <= 35'd34288443811;
	bram[43] <= 35'd34285011373;
	bram[44] <= 35'd34281497015;
	bram[45] <= 35'd34277900737;
	bram[46] <= 35'd34274222538;
	bram[47] <= 35'd34270470613;
	bram[48] <= 35'd34266628574;
	bram[49] <= 35'd34262712808;
	bram[50] <= 35'd34258715122;
	bram[51] <= 35'd34254635516;
	bram[52] <= 35'd34250473989;
	bram[53] <= 35'd34246238736;
	bram[54] <= 35'd34241913369;
	bram[55] <= 35'd34237514275;
	bram[56] <= 35'd34233033261;
	bram[57] <= 35'd34228470327;
	bram[58] <= 35'd34223825472;
	bram[59] <= 35'd34219106891;
	bram[60] <= 35'd34214298196;
	bram[61] <= 35'd34209415774;
	bram[62] <= 35'd34204451432;
	bram[63] <= 35'd34199405170;
	bram[64] <= 35'd34194276987;
	bram[65] <= 35'd34189075078;
	bram[66] <= 35'd34183783055;
	bram[67] <= 35'd34178417305;
	bram[68] <= 35'd34172969635;
	bram[69] <= 35'd34167440044;
	bram[70] <= 35'd34161836727;
	bram[71] <= 35'd34156143296;
	bram[72] <= 35'd34150376138;
	bram[73] <= 35'd34144527060;
	bram[74] <= 35'd34138596062;
	bram[75] <= 35'd34132583143;
	bram[76] <= 35'd34126496497;
	bram[77] <= 35'd34120327932;
	bram[78] <= 35'd34114069252;
	bram[79] <= 35'd34107745039;
	bram[80] <= 35'd34101330713;
	bram[81] <= 35'd34094834466;
	bram[82] <= 35'd34088264492;
	bram[83] <= 35'd34081612598;
	bram[84] <= 35'd34074878783;
	bram[85] <= 35'd34068071242;
	bram[86] <= 35'd34061173587;
	bram[87] <= 35'd34054202205;
	bram[88] <= 35'd34047148903;
	bram[89] <= 35'd34040013680;
	bram[90] <= 35'd34032804731;
	bram[91] <= 35'd34025505668;
	bram[92] <= 35'd34018132878;
	bram[93] <= 35'd34010678167;
	bram[94] <= 35'd34003149730;
	bram[95] <= 35'd33995531179;
	bram[96] <= 35'd33987838901;
	bram[97] <= 35'd33980064703;
	bram[98] <= 35'd33972208584;
	bram[99] <= 35'd33964278738;
	bram[100] <= 35'd33956266972;
	bram[101] <= 35'd33948173286;
	bram[102] <= 35'd33939997679;
	bram[103] <= 35'd33931748346;
	bram[104] <= 35'd33923408899;
	bram[105] <= 35'd33914995724;
	bram[106] <= 35'd33906508823;
	bram[107] <= 35'd33897931808;
	bram[108] <= 35'd33889281066;
	bram[109] <= 35'd33880548404;
	bram[110] <= 35'd33871733821;
	bram[111] <= 35'd33862845511;
	bram[112] <= 35'd33853875281;
	bram[113] <= 35'd33844823130;
	bram[114] <= 35'd33835697253;
	bram[115] <= 35'd33826481262;
	bram[116] <= 35'd33817191543;
	bram[117] <= 35'd33807828098;
	bram[118] <= 35'd33798374539;
	bram[119] <= 35'd33788847253;
	bram[120] <= 35'd33779238046;
	bram[121] <= 35'd33769555112;
	bram[122] <= 35'd33759790258;
	bram[123] <= 35'd33749943484;
	bram[124] <= 35'd33740014789;
	bram[125] <= 35'd33730012367;
	bram[126] <= 35'd33719928025;
	bram[127] <= 35'd33709761762;
	bram[128] <= 35'd33699521772;
	bram[129] <= 35'd33689199862;
	bram[130] <= 35'd33678796032;
	bram[131] <= 35'd33668310281;
	bram[132] <= 35'd33657750802;
	bram[133] <= 35'd33647117597;
	bram[134] <= 35'd33636394278;
	bram[135] <= 35'd33625597232;
	bram[136] <= 35'd33614718265;
	bram[137] <= 35'd33603765571;
	bram[138] <= 35'd33592730957;
	bram[139] <= 35'd33581614422;
	bram[140] <= 35'd33570424160;
	bram[141] <= 35'd33559151978;
	bram[142] <= 35'd33547797875;
	bram[143] <= 35'd33536370045;
	bram[144] <= 35'd33524860294;
	bram[145] <= 35'd33513276816;
	bram[146] <= 35'd33501611418;
	bram[147] <= 35'd33489864099;
	bram[148] <= 35'd33478043053;
	bram[149] <= 35'd33466140087;
	bram[150] <= 35'd33454155200;
	bram[151] <= 35'd33442096586;
	bram[152] <= 35'd33429956051;
	bram[153] <= 35'd33417741789;
	bram[154] <= 35'd33405445607;
	bram[155] <= 35'd33393067504;
	bram[156] <= 35'd33380615674;
	bram[157] <= 35'd33368081923;
	bram[158] <= 35'd33355474445;
	bram[159] <= 35'd33342785047;
	bram[160] <= 35'd33330013728;
	bram[161] <= 35'd33317168682;
	bram[162] <= 35'd33304241715;
	bram[163] <= 35'd33291241021;
	bram[164] <= 35'd33278158406;
	bram[165] <= 35'd33265002064;
	bram[166] <= 35'd33251763802;
	bram[167] <= 35'd33238443619;
	bram[168] <= 35'd33225049708;
	bram[169] <= 35'd33211582070;
	bram[170] <= 35'd33198032512;
	bram[171] <= 35'd33184401033;
	bram[172] <= 35'd33170695827;
	bram[173] <= 35'd33156908700;
	bram[174] <= 35'd33143047846;
	bram[175] <= 35'd33129105071;
	bram[176] <= 35'd33115088569;
	bram[177] <= 35'd33100990146;
	bram[178] <= 35'd33086817996;
	bram[179] <= 35'd33072563925;
	bram[180] <= 35'd33058236127;
	bram[181] <= 35'd33043826408;
	bram[182] <= 35'd33029342962;
	bram[183] <= 35'd33014777595;
	bram[184] <= 35'd33000138501;
	bram[185] <= 35'd32985417486;
	bram[186] <= 35'd32970622744;
	bram[187] <= 35'd32955746081;
	bram[188] <= 35'd32940795691;
	bram[189] <= 35'd32925763380;
	bram[190] <= 35'd32910657341;
	bram[191] <= 35'd32895477575;
	bram[192] <= 35'd32880215889;
	bram[193] <= 35'd32864872282;
	bram[194] <= 35'd32849454947;
	bram[195] <= 35'd32833963885;
	bram[196] <= 35'd32818390902;
	bram[197] <= 35'd32802744191;
	bram[198] <= 35'd32787023753;
	bram[199] <= 35'd32771221395;
	bram[200] <= 35'd32755337115;
	bram[201] <= 35'd32739387302;
	bram[202] <= 35'd32723347374;
	bram[203] <= 35'd32707241912;
	bram[204] <= 35'd32691054530;
	bram[205] <= 35'd32674785226;
	bram[206] <= 35'd32658450389;
	bram[207] <= 35'd32642025437;
	bram[208] <= 35'd32625534951;
	bram[209] <= 35'd32608962544;
	bram[210] <= 35'd32592316410;
	bram[211] <= 35'd32575588355;
	bram[212] <= 35'd32558786572;
	bram[213] <= 35'd32541911062;
	bram[214] <= 35'd32524953631;
	bram[215] <= 35'd32507922472;
	bram[216] <= 35'd32490817586;
	bram[217] <= 35'd32473630779;
	bram[218] <= 35'd32456370244;
	bram[219] <= 35'd32439035982;
	bram[220] <= 35'd32421619799;
	bram[221] <= 35'd32404129888;
	bram[222] <= 35'd32386566250;
	bram[223] <= 35'd32368920691;
	bram[224] <= 35'd32351201404;
	bram[225] <= 35'd32333408390;
	bram[226] <= 35'd32315533454;
	bram[227] <= 35'd32297592984;
	bram[228] <= 35'd32279570594;
	bram[229] <= 35'd32261466282;
	bram[230] <= 35'd32243296436;
	bram[231] <= 35'd32225044669;
	bram[232] <= 35'd32206719175;
	bram[233] <= 35'd32188311759;
	bram[234] <= 35'd32169838809;
	bram[235] <= 35'd32151283938;
	bram[236] <= 35'd32132655339;
	bram[237] <= 35'd32113953013;
	bram[238] <= 35'd32095168766;
	bram[239] <= 35'd32076310791;
	bram[240] <= 35'd32057379088;
	bram[241] <= 35'd32038373657;
	bram[242] <= 35'd32019294499;
	bram[243] <= 35'd32000133419;
	bram[244] <= 35'd31980906805;
	bram[245] <= 35'd31961598270;
	bram[246] <= 35'd31942216008;
	bram[247] <= 35'd31922751824;
	bram[248] <= 35'd31903222106;
	bram[249] <= 35'd31883610467;
	bram[250] <= 35'd31863925100;
	bram[251] <= 35'd31844166005;
	bram[252] <= 35'd31824333182;
	bram[253] <= 35'd31804426631;
	bram[254] <= 35'd31784446353;
	bram[255] <= 35'd31764384153;
	bram[256] <= 35'd31744256419;
	bram[257] <= 35'd31724046764;
	bram[258] <= 35'd31703763381;
	bram[259] <= 35'd31683406270;
	bram[260] <= 35'd31662975431;
	bram[261] <= 35'd31642470864;
	bram[262] <= 35'd31621892570;
	bram[263] <= 35'd31601232354;
	bram[264] <= 35'd31580506603;
	bram[265] <= 35'd31559707125;
	bram[266] <= 35'd31538825726;
	bram[267] <= 35'd31517870598;
	bram[268] <= 35'd31496849936;
	bram[269] <= 35'd31475747353;
	bram[270] <= 35'd31454571041;
	bram[271] <= 35'd31433329195;
	bram[272] <= 35'd31412005428;
	bram[273] <= 35'd31390607933;
	bram[274] <= 35'd31369136710;
	bram[275] <= 35'd31347591759;
	bram[276] <= 35'd31325973080;
	bram[277] <= 35'd31304280672;
	bram[278] <= 35'd31282522730;
	bram[279] <= 35'd31260682867;
	bram[280] <= 35'd31238769276;
	bram[281] <= 35'd31216781957;
	bram[282] <= 35'd31194720909;
	bram[283] <= 35'd31172594327;
	bram[284] <= 35'd31150385824;
	bram[285] <= 35'd31128103592;
	bram[286] <= 35'd31105755826;
	bram[287] <= 35'd31083326138;
	bram[288] <= 35'd31060830915;
	bram[289] <= 35'd31038261965;
	bram[290] <= 35'd31015611093;
	bram[291] <= 35'd30992894686;
	bram[292] <= 35'd30970104551;
	bram[293] <= 35'd30947240688;
	bram[294] <= 35'd30924303096;
	bram[295] <= 35'd30901299970;
	bram[296] <= 35'd30878214922;
	bram[297] <= 35'd30855064340;
	bram[298] <= 35'd30831831836;
	bram[299] <= 35'd30808533797;
	bram[300] <= 35'd30785162030;
	bram[301] <= 35'd30761716535;
	bram[302] <= 35'd30738197311;
	bram[303] <= 35'd30714612553;
	bram[304] <= 35'd30690945873;
	bram[305] <= 35'd30667213658;
	bram[306] <= 35'd30643407715;
	bram[307] <= 35'd30619528043;
	bram[308] <= 35'd30595582837;
	bram[309] <= 35'd30571555709;
	bram[310] <= 35'd30547463046;
	bram[311] <= 35'd30523296654;
	bram[312] <= 35'd30499064728;
	bram[313] <= 35'd30474750880;
	bram[314] <= 35'd30450371497;
	bram[315] <= 35'd30425918386;
	bram[316] <= 35'd30401391546;
	bram[317] <= 35'd30376799171;
	bram[318] <= 35'd30352133068;
	bram[319] <= 35'd30327393237;
	bram[320] <= 35'd30302579677;
	bram[321] <= 35'd30277700582;
	bram[322] <= 35'd30252747759;
	bram[323] <= 35'd30227721207;
	bram[324] <= 35'd30202629120;
	bram[325] <= 35'd30177463305;
	bram[326] <= 35'd30152223762;
	bram[327] <= 35'd30126910490;
	bram[328] <= 35'd30101531682;
	bram[329] <= 35'd30076087340;
	bram[330] <= 35'd30050561076;
	bram[331] <= 35'd30024969276;
	bram[332] <= 35'd29999311941;
	bram[333] <= 35'd29973580878;
	bram[334] <= 35'd29947776087;
	bram[335] <= 35'd29921897567;
	bram[336] <= 35'd29895953511;
	bram[337] <= 35'd29869943920;
	bram[338] <= 35'd29843860601;
	bram[339] <= 35'd29817703553;
	bram[340] <= 35'd29791480970;
	bram[341] <= 35'd29765184659;
	bram[342] <= 35'd29738814619;
	bram[343] <= 35'd29712379043;
	bram[344] <= 35'd29685877932;
	bram[345] <= 35'd29659303093;
	bram[346] <= 35'd29632654525;
	bram[347] <= 35'd29605940421;
	bram[348] <= 35'd29579160782;
	bram[349] <= 35'd29552307415;
	bram[350] <= 35'd29525380319;
	bram[351] <= 35'd29498387687;
	bram[352] <= 35'd29471329520;
	bram[353] <= 35'd29444197625;
	bram[354] <= 35'd29416992001;
	bram[355] <= 35'd29389720841;
	bram[356] <= 35'd29362384146;
	bram[357] <= 35'd29334973722;
	bram[358] <= 35'd29307497762;
	bram[359] <= 35'd29279956267;
	bram[360] <= 35'd29252341044;
	bram[361] <= 35'd29224652092;
	bram[362] <= 35'd29196897604;
	bram[363] <= 35'd29169077580;
	bram[364] <= 35'd29141192021;
	bram[365] <= 35'd29113232734;
	bram[366] <= 35'd29085199717;
	bram[367] <= 35'd29057109358;
	bram[368] <= 35'd29028945270;
	bram[369] <= 35'd29000715647;
	bram[370] <= 35'd28972412295;
	bram[371] <= 35'd28944043407;
	bram[372] <= 35'd28915608984;
	bram[373] <= 35'd28887100832;
	bram[374] <= 35'd28858527144;
	bram[375] <= 35'd28829887921;
	bram[376] <= 35'd28801174968;
	bram[377] <= 35'd28772404673;
	bram[378] <= 35'd28743560650;
	bram[379] <= 35'd28714642897;
	bram[380] <= 35'd28685667802;
	bram[381] <= 35'd28656618978;
	bram[382] <= 35'd28627504618;
	bram[383] <= 35'd28598324723;
	bram[384] <= 35'd28569071098;
	bram[385] <= 35'd28539760131;
	bram[386] <= 35'd28510375435;
	bram[387] <= 35'd28480925203;
	bram[388] <= 35'd28451409436;
	bram[389] <= 35'd28421819939;
	bram[390] <= 35'd28392173100;
	bram[391] <= 35'd28362452532;
	bram[392] <= 35'd28332666428;
	bram[393] <= 35'd28302814788;
	bram[394] <= 35'd28272897612;
	bram[395] <= 35'd28242914900;
	bram[396] <= 35'd28212866653;
	bram[397] <= 35'd28182744676;
	bram[398] <= 35'd28152565357;
	bram[399] <= 35'd28122312309;
	bram[400] <= 35'd28091993724;
	bram[401] <= 35'd28061617797;
	bram[402] <= 35'd28031168141;
	bram[403] <= 35'd28000652949;
	bram[404] <= 35'd27970072221;
	bram[405] <= 35'd27939425957;
	bram[406] <= 35'd27908714157;
	bram[407] <= 35'd27877936821;
	bram[408] <= 35'd27847093949;
	bram[409] <= 35'd27816185541;
	bram[410] <= 35'd27785211597;
	bram[411] <= 35'd27754172117;
	bram[412] <= 35'd27723067101;
	bram[413] <= 35'd27691896549;
	bram[414] <= 35'd27660660460;
	bram[415] <= 35'd27629367029;
	bram[416] <= 35'd27597999869;
	bram[417] <= 35'd27566567173;
	bram[418] <= 35'd27535068940;
	bram[419] <= 35'd27503513364;
	bram[420] <= 35'd27471892253;
	bram[421] <= 35'd27440197412;
	bram[422] <= 35'd27408445228;
	bram[423] <= 35'd27376627508;
	bram[424] <= 35'd27344744252;
	bram[425] <= 35'd27312795459;
	bram[426] <= 35'd27280789324;
	bram[427] <= 35'd27248709459;
	bram[428] <= 35'd27216572251;
	bram[429] <= 35'd27184369507;
	bram[430] <= 35'd27152101227;
	bram[431] <= 35'd27119767410;
	bram[432] <= 35'd27087376250;
	bram[433] <= 35'd27054919555;
	bram[434] <= 35'd27022389129;
	bram[435] <= 35'd26989809554;
	bram[436] <= 35'd26957156249;
	bram[437] <= 35'd26924445601;
	bram[438] <= 35'd26891669417;
	bram[439] <= 35'd26858827696;
	bram[440] <= 35'd26825928633;
	bram[441] <= 35'd26792955840;
	bram[442] <= 35'd26759925703;
	bram[443] <= 35'd26726838223;
	bram[444] <= 35'd26693685207;
	bram[445] <= 35'd26660466655;
	bram[446] <= 35'd26627182566;
	bram[447] <= 35'd26593841134;
	bram[448] <= 35'd26560434165;
	bram[449] <= 35'd26526969854;
	bram[450] <= 35'd26493431812;
	bram[451] <= 35'd26459844621;
	bram[452] <= 35'd26426183699;
	bram[453] <= 35'd26392473628;
	bram[454] <= 35'd26358689827;
	bram[455] <= 35'd26324848683;
	bram[456] <= 35'd26290942002;
	bram[457] <= 35'd26256977978;
	bram[458] <= 35'd26222948417;
	bram[459] <= 35'd26188861513;
	bram[460] <= 35'd26154709072;
	bram[461] <= 35'd26120499288;
	bram[462] <= 35'd26086223967;
	bram[463] <= 35'd26051891303;
	bram[464] <= 35'd26017493102;
	bram[465] <= 35'd25983037558;
	bram[466] <= 35'd25948516477;
	bram[467] <= 35'd25913938052;
	bram[468] <= 35'd25879302284;
	bram[469] <= 35'd25844600980;
	bram[470] <= 35'd25809834139;
	bram[471] <= 35'd25775009954;
	bram[472] <= 35'd25740128426;
	bram[473] <= 35'd25705181361;
	bram[474] <= 35'd25670176952;
	bram[475] <= 35'd25635115200;
	bram[476] <= 35'd25599987911;
	bram[477] <= 35'd25564803279;
	bram[478] <= 35'd25529553109;
	bram[479] <= 35'd25494253789;
	bram[480] <= 35'd25458888933;
	bram[481] <= 35'd25423458540;
	bram[482] <= 35'd25387970803;
	bram[483] <= 35'd25352425722;
	bram[484] <= 35'd25316823298;
	bram[485] <= 35'd25281155337;
	bram[486] <= 35'd25245430032;
	bram[487] <= 35'd25209647383;
	bram[488] <= 35'd25173807391;
	bram[489] <= 35'd25137901861;
	bram[490] <= 35'd25101947181;
	bram[491] <= 35'd25065926965;
	bram[492] <= 35'd25029841211;
	bram[493] <= 35'd24993706307;
	bram[494] <= 35'd24957505865;
	bram[495] <= 35'd24921256273;
	bram[496] <= 35'd24884941144;
	bram[497] <= 35'd24848568672;
	bram[498] <= 35'd24812130662;
	bram[499] <= 35'd24775643501;
	bram[500] <= 35'd24739098997;
	bram[501] <= 35'd24702488956;
	bram[502] <= 35'd24665821570;
	bram[503] <= 35'd24629105034;
	bram[504] <= 35'd24592322961;
	bram[505] <= 35'd24555483544;
	bram[506] <= 35'd24518586783;
	bram[507] <= 35'd24481632678;
	bram[508] <= 35'd24444621229;
	bram[509] <= 35'd24407552436;
	bram[510] <= 35'd24370426299;
	bram[511] <= 35'd24333242818;
	bram[512] <= 35'd24296001993;
	bram[513] <= 35'd24258703824;
	bram[514] <= 35'd24221348311;
	bram[515] <= 35'd24183935454;
	bram[516] <= 35'd24146465252;
	bram[517] <= 35'd24108945900;
	bram[518] <= 35'd24071361011;
	bram[519] <= 35'd24033718777;
	bram[520] <= 35'd23996027393;
	bram[521] <= 35'd23958270471;
	bram[522] <= 35'd23920464398;
	bram[523] <= 35'd23882600981;
	bram[524] <= 35'd23844680220;
	bram[525] <= 35'd23806702115;
	bram[526] <= 35'd23768666666;
	bram[527] <= 35'd23730573872;
	bram[528] <= 35'd23692431927;
	bram[529] <= 35'd23654232638;
	bram[530] <= 35'd23615976005;
	bram[531] <= 35'd23577662028;
	bram[532] <= 35'd23539290706;
	bram[533] <= 35'd23500870233;
	bram[534] <= 35'd23462392416;
	bram[535] <= 35'd23423857254;
	bram[536] <= 35'd23385272941;
	bram[537] <= 35'd23346631284;
	bram[538] <= 35'd23307932283;
	bram[539] <= 35'd23269175937;
	bram[540] <= 35'd23230370440;
	bram[541] <= 35'd23191507599;
	bram[542] <= 35'd23152587413;
	bram[543] <= 35'd23113618076;
	bram[544] <= 35'd23074591395;
	bram[545] <= 35'd23035507369;
	bram[546] <= 35'd22996374192;
	bram[547] <= 35'd22957183670;
	bram[548] <= 35'd22917943997;
	bram[549] <= 35'd22878646980;
	bram[550] <= 35'd22839292618;
	bram[551] <= 35'd22799889105;
	bram[552] <= 35'd22760428247;
	bram[553] <= 35'd22720918237;
	bram[554] <= 35'd22681359077;
	bram[555] <= 35'd22641734378;
	bram[556] <= 35'd22602068722;
	bram[557] <= 35'd22562337527;
	bram[558] <= 35'd22522565375;
	bram[559] <= 35'd22482727684;
	bram[560] <= 35'd22442849035;
	bram[561] <= 35'd22402913042;
	bram[562] <= 35'd22362919704;
	bram[563] <= 35'd22322877214;
	bram[564] <= 35'd22282785573;
	bram[565] <= 35'd22242636587;
	bram[566] <= 35'd22202438450;
	bram[567] <= 35'd22162182967;
	bram[568] <= 35'd22121886527;
	bram[569] <= 35'd22081524548;
	bram[570] <= 35'd22041121611;
	bram[571] <= 35'd22000661329;
	bram[572] <= 35'd21960151896;
	bram[573] <= 35'd21919585118;
	bram[574] <= 35'd21878969188;
	bram[575] <= 35'd21838304106;
	bram[576] <= 35'd21797589873;
	bram[577] <= 35'd21756818295;
	bram[578] <= 35'd21715997565;
	bram[579] <= 35'd21675127683;
	bram[580] <= 35'd21634208650;
	bram[581] <= 35'd21593232272;
	bram[582] <= 35'd21552206742;
	bram[583] <= 35'd21511132060;
	bram[584] <= 35'd21470008226;
	bram[585] <= 35'd21428835241;
	bram[586] <= 35'd21387604910;
	bram[587] <= 35'd21346333621;
	bram[588] <= 35'd21305004987;
	bram[589] <= 35'd21263627201;
	bram[590] <= 35'd21222200263;
	bram[591] <= 35'd21180724173;
	bram[592] <= 35'd21139198932;
	bram[593] <= 35'd21097616345;
	bram[594] <= 35'd21055992799;
	bram[595] <= 35'd21014320102;
	bram[596] <= 35'd20972590059;
	bram[597] <= 35'd20930819057;
	bram[598] <= 35'd20888998904;
	bram[599] <= 35'd20847121405;
	bram[600] <= 35'd20805202948;
	bram[601] <= 35'd20763227145;
	bram[602] <= 35'd20721210383;
	bram[603] <= 35'd20679144469;
	bram[604] <= 35'd20637029404;
	bram[605] <= 35'd20594856993;
	bram[606] <= 35'd20552643623;
	bram[607] <= 35'd20510381101;
	bram[608] <= 35'd20468069426;
	bram[609] <= 35'd20425716793;
	bram[610] <= 35'd20383306814;
	bram[611] <= 35'd20340855877;
	bram[612] <= 35'd20298347594;
	bram[613] <= 35'd20255798352;
	bram[614] <= 35'd20213199958;
	bram[615] <= 35'd20170552411;
	bram[616] <= 35'd20127863906;
	bram[617] <= 35'd20085118055;
	bram[618] <= 35'd20042331245;
	bram[619] <= 35'd19999495282;
	bram[620] <= 35'd19956618361;
	bram[621] <= 35'd19913684094;
	bram[622] <= 35'd19870708867;
	bram[623] <= 35'd19827692682;
	bram[624] <= 35'd19784619151;
	bram[625] <= 35'd19741504661;
	bram[626] <= 35'd19698341018;
	bram[627] <= 35'd19655136417;
	bram[628] <= 35'd19611874469;
	bram[629] <= 35'd19568579756;
	bram[630] <= 35'd19525227697;
	bram[631] <= 35'd19481834678;
	bram[632] <= 35'd19438400701;
	bram[633] <= 35'd19394909377;
	bram[634] <= 35'd19351385288;
	bram[635] <= 35'd19307803852;
	bram[636] <= 35'd19264189651;
	bram[637] <= 35'd19220518104;
	bram[638] <= 35'd19176805597;
	bram[639] <= 35'd19133052131;
	bram[640] <= 35'd19089249513;
	bram[641] <= 35'd19045397741;
	bram[642] <= 35'd19001513204;
	bram[643] <= 35'd18957571320;
	bram[644] <= 35'd18913596671;
	bram[645] <= 35'd18869564675;
	bram[646] <= 35'd18825499913;
	bram[647] <= 35'd18781385999;
	bram[648] <= 35'd18737222932;
	bram[649] <= 35'd18693018905;
	bram[650] <= 35'd18648773918;
	bram[651] <= 35'd18604487972;
	bram[652] <= 35'd18560152873;
	bram[653] <= 35'd18515776815;
	bram[654] <= 35'd18471351604;
	bram[655] <= 35'd18426885433;
	bram[656] <= 35'd18382378302;
	bram[657] <= 35'd18337830212;
	bram[658] <= 35'd18293232969;
	bram[659] <= 35'd18248594766;
	bram[660] <= 35'd18203915603;
	bram[661] <= 35'd18159195481;
	bram[662] <= 35'd18114426206;
	bram[663] <= 35'd18069615971;
	bram[664] <= 35'd18024764776;
	bram[665] <= 35'd17979872621;
	bram[666] <= 35'd17934939507;
	bram[667] <= 35'd17889957240;
	bram[668] <= 35'd17844934012;
	bram[669] <= 35'd17799878018;
	bram[670] <= 35'd17754772871;
	bram[671] <= 35'd17709626764;
	bram[672] <= 35'd17664439697;
	bram[673] <= 35'd17619211671;
	bram[674] <= 35'd17573934491;
	bram[675] <= 35'd17528624544;
	bram[676] <= 35'd17483273638;
	bram[677] <= 35'd17437873578;
	bram[678] <= 35'd17392440751;
	bram[679] <= 35'd17346966964;
	bram[680] <= 35'd17301452218;
	bram[681] <= 35'd17255888318;
	bram[682] <= 35'd17210291651;
	bram[683] <= 35'd17164654024;
	bram[684] <= 35'd17118975437;
	bram[685] <= 35'd17073255890;
	bram[686] <= 35'd17027495383;
	bram[687] <= 35'd16981693916;
	bram[688] <= 35'd16935851488;
	bram[689] <= 35'd16889976294;
	bram[690] <= 35'd16844051946;
	bram[691] <= 35'd16798094831;
	bram[692] <= 35'd16752096756;
	bram[693] <= 35'd16706057720;
	bram[694] <= 35'd16659985918;
	bram[695] <= 35'd16613864962;
	bram[696] <= 35'd16567711239;
	bram[697] <= 35'd16521516556;
	bram[698] <= 35'd16475280912;
	bram[699] <= 35'd16429012502;
	bram[700] <= 35'd16382694937;
	bram[701] <= 35'd16336352799;
	bram[702] <= 35'd16289961507;
	bram[703] <= 35'd16243537448;
	bram[704] <= 35'd16197072429;
	bram[705] <= 35'd16150566449;
	bram[706] <= 35'd16104027702;
	bram[707] <= 35'd16057447994;
	bram[708] <= 35'd16010835519;
	bram[709] <= 35'd15964182084;
	bram[710] <= 35'd15917487688;
	bram[711] <= 35'd15870760525;
	bram[712] <= 35'd15823992401;
	bram[713] <= 35'd15777191510;
	bram[714] <= 35'd15730349659;
	bram[715] <= 35'd15683466847;
	bram[716] <= 35'd15636551267;
	bram[717] <= 35'd15589602920;
	bram[718] <= 35'd15542613612;
	bram[719] <= 35'd15495591537;
	bram[720] <= 35'd15448528501;
	bram[721] <= 35'd15401432698;
	bram[722] <= 35'd15354295934;
	bram[723] <= 35'd15307126402;
	bram[724] <= 35'd15259924103;
	bram[725] <= 35'd15212680843;
	bram[726] <= 35'd15165404816;
	bram[727] <= 35'd15118087828;
	bram[728] <= 35'd15070738072;
	bram[729] <= 35'd15023355548;
	bram[730] <= 35'd14975940257;
	bram[731] <= 35'd14928484005;
	bram[732] <= 35'd14880994986;
	bram[733] <= 35'd14833465005;
	bram[734] <= 35'd14785910450;
	bram[735] <= 35'd14738314934;
	bram[736] <= 35'd14690686651;
	bram[737] <= 35'd14643017406;
	bram[738] <= 35'd14595323587;
	bram[739] <= 35'd14547588807;
	bram[740] <= 35'd14499821259;
	bram[741] <= 35'd14452020943;
	bram[742] <= 35'd14404187860;
	bram[743] <= 35'd14356313815;
	bram[744] <= 35'd14308415196;
	bram[745] <= 35'd14260475616;
	bram[746] <= 35'd14212503267;
	bram[747] <= 35'd14164506344;
	bram[748] <= 35'd14116468460;
	bram[749] <= 35'd14068397808;
	bram[750] <= 35'd14020294388;
	bram[751] <= 35'd13972158200;
	bram[752] <= 35'd13923989244;
	bram[753] <= 35'd13875787520;
	bram[754] <= 35'd13827553028;
	bram[755] <= 35'd13779285768;
	bram[756] <= 35'd13730985740;
	bram[757] <= 35'd13682652944;
	bram[758] <= 35'd13634287379;
	bram[759] <= 35'd13585897240;
	bram[760] <= 35'd13537466140;
	bram[761] <= 35'd13489002271;
	bram[762] <= 35'd13440513827;
	bram[763] <= 35'd13391992615;
	bram[764] <= 35'd13343438635;
	bram[765] <= 35'd13294851887;
	bram[766] <= 35'd13246232370;
	bram[767] <= 35'd13197588279;
	bram[768] <= 35'd13148903226;
	bram[769] <= 35'd13100193598;
	bram[770] <= 35'd13051451201;
	bram[771] <= 35'd13002684230;
	bram[772] <= 35'd12953876297;
	bram[773] <= 35'd12905043789;
	bram[774] <= 35'd12856178512;
	bram[775] <= 35'd12807288660;
	bram[776] <= 35'd12758366040;
	bram[777] <= 35'd12709410651;
	bram[778] <= 35'd12660430688;
	bram[779] <= 35'd12611409762;
	bram[780] <= 35'd12562372455;
	bram[781] <= 35'd12513294186;
	bram[782] <= 35'd12464191341;
	bram[783] <= 35'd12415063921;
	bram[784] <= 35'd12365903733;
	bram[785] <= 35'd12316710776;
	bram[786] <= 35'd12267493244;
	bram[787] <= 35'd12218242943;
	bram[788] <= 35'd12168968067;
	bram[789] <= 35'd12119660422;
	bram[790] <= 35'd12070328201;
	bram[791] <= 35'd12020971405;
	bram[792] <= 35'd11971581841;
	bram[793] <= 35'd11922159508;
	bram[794] <= 35'd11872712599;
	bram[795] <= 35'd11823241115;
	bram[796] <= 35'd11773736862;
	bram[797] <= 35'd11724208034;
	bram[798] <= 35'd11674646437;
	bram[799] <= 35'd11625060264;
	bram[800] <= 35'd11575449515;
	bram[801] <= 35'd11525814191;
	bram[802] <= 35'd11476146098;
	bram[803] <= 35'd11426453430;
	bram[804] <= 35'd11376727993;
	bram[805] <= 35'd11326977979;
	bram[806] <= 35'd11277211584;
	bram[807] <= 35'd11227404226;
	bram[808] <= 35'd11177580486;
	bram[809] <= 35'd11127723977;
	bram[810] <= 35'd11077842892;
	bram[811] <= 35'd11027937231;
	bram[812] <= 35'd10978006994;
	bram[813] <= 35'd10928052181;
	bram[814] <= 35'd10878072793;
	bram[815] <= 35'd10828060636;
	bram[816] <= 35'd10778023903;
	bram[817] <= 35'd10727962593;
	bram[818] <= 35'd10677884901;
	bram[819] <= 35'd10627774440;
	bram[820] <= 35'd10577639403;
	bram[821] <= 35'd10527479790;
	bram[822] <= 35'd10477295601;
	bram[823] <= 35'd10427086837;
	bram[824] <= 35'd10376845303;
	bram[825] <= 35'd10326587386;
	bram[826] <= 35'd10276304893;
	bram[827] <= 35'd10225997823;
	bram[828] <= 35'd10175674371;
	bram[829] <= 35'd10125318150;
	bram[830] <= 35'd10074937353;
	bram[831] <= 35'd10024531979;
	bram[832] <= 35'd9974110222;
	bram[833] <= 35'd9923663890;
	bram[834] <= 35'd9873184788;
	bram[835] <= 35'd9822689303;
	bram[836] <= 35'd9772169241;
	bram[837] <= 35'd9721632797;
	bram[838] <= 35'd9671063583;
	bram[839] <= 35'd9620477986;
	bram[840] <= 35'd9569867813;
	bram[841] <= 35'd9519233063;
	bram[842] <= 35'd9468581931;
	bram[843] <= 35'd9417898028;
	bram[844] <= 35'd9367205936;
	bram[845] <= 35'd9316481074;
	bram[846] <= 35'd9265739829;
	bram[847] <= 35'd9214974008;
	bram[848] <= 35'd9164183610;
	bram[849] <= 35'd9113376829;
	bram[850] <= 35'd9062545471;
	bram[851] <= 35'd9011697730;
	bram[852] <= 35'd8960825413;
	bram[853] <= 35'd8909928519;
	bram[854] <= 35'd8859015242;
	bram[855] <= 35'd8808077388;
	bram[856] <= 35'd8757123151;
	bram[857] <= 35'd8706144337;
	bram[858] <= 35'd8655149140;
	bram[859] <= 35'd8604129366;
	bram[860] <= 35'd8553093209;
	bram[861] <= 35'd8502032475;
	bram[862] <= 35'd8450955358;
	bram[863] <= 35'd8399853664;
	bram[864] <= 35'd8348735586;
	bram[865] <= 35'd8297601125;
	bram[866] <= 35'd8246442087;
	bram[867] <= 35'd8195266665;
	bram[868] <= 35'd8144074860;
	bram[869] <= 35'd8092858478;
	bram[870] <= 35'd8041625713;
	bram[871] <= 35'd7990368370;
	bram[872] <= 35'd7939102837;
	bram[873] <= 35'd7887812728;
	bram[874] <= 35'd7836498041;
	bram[875] <= 35'd7785175164;
	bram[876] <= 35'd7733827710;
	bram[877] <= 35'd7682463872;
	bram[878] <= 35'd7631083650;
	bram[879] <= 35'd7579687045;
	bram[880] <= 35'd7528265863;
	bram[881] <= 35'd7476828297;
	bram[882] <= 35'd7425374347;
	bram[883] <= 35'd7373904013;
	bram[884] <= 35'd7322417295;
	bram[885] <= 35'd7270914193;
	bram[886] <= 35'd7219394708;
	bram[887] <= 35'd7167850645;
	bram[888] <= 35'd7116298392;
	bram[889] <= 35'd7064721561;
	bram[890] <= 35'd7013136540;
	bram[891] <= 35'd6961526941;
	bram[892] <= 35'd6909909152;
	bram[893] <= 35'd6858266785;
	bram[894] <= 35'd6806616228;
	bram[895] <= 35'd6754941093;
	bram[896] <= 35'd6703257767;
	bram[897] <= 35'd6651558058;
	bram[898] <= 35'd6599833771;
	bram[899] <= 35'd6548101293;
	bram[900] <= 35'd6496352431;
	bram[901] <= 35'd6444587184;
	bram[902] <= 35'd6392813747;
	bram[903] <= 35'd6341015732;
	bram[904] <= 35'd6289209526;
	bram[905] <= 35'd6237386936;
	bram[906] <= 35'd6185547962;
	bram[907] <= 35'd6133692604;
	bram[908] <= 35'd6081820861;
	bram[909] <= 35'd6029940927;
	bram[910] <= 35'd5978044609;
	bram[911] <= 35'd5926131906;
	bram[912] <= 35'd5874211012;
	bram[913] <= 35'd5822273734;
	bram[914] <= 35'd5770320071;
	bram[915] <= 35'd5718358217;
	bram[916] <= 35'd5666379979;
	bram[917] <= 35'd5614385356;
	bram[918] <= 35'd5562382542;
	bram[919] <= 35'd5510363344;
	bram[920] <= 35'd5458327761;
	bram[921] <= 35'd5406283986;
	bram[922] <= 35'd5354232021;
	bram[923] <= 35'd5302155477;
	bram[924] <= 35'd5250078935;
	bram[925] <= 35'd5197986009;
	bram[926] <= 35'd5145876698;
	bram[927] <= 35'd5093759196;
	bram[928] <= 35'd5041625309;
	bram[929] <= 35'd4989483230;
	bram[930] <= 35'd4937332960;
	bram[931] <= 35'd4885166306;
	bram[932] <= 35'd4832983266;
	bram[933] <= 35'd4780800229;
	bram[934] <= 35'd4728592613;
	bram[935] <= 35'd4676384999;
	bram[936] <= 35'd4624161000;
	bram[937] <= 35'd4571928809;
	bram[938] <= 35'd4519688427;
	bram[939] <= 35'd4467431660;
	bram[940] <= 35'd4415166701;
	bram[941] <= 35'd4362893551;
	bram[942] <= 35'd4310604016;
	bram[943] <= 35'd4258306289;
	bram[944] <= 35'd4206000370;
	bram[945] <= 35'd4153686259;
	bram[946] <= 35'd4101363957;
	bram[947] <= 35'd4049025269;
	bram[948] <= 35'd3996686583;
	bram[949] <= 35'd3944331512;
	bram[950] <= 35'd3891968249;
	bram[951] <= 35'd3839596795;
	bram[952] <= 35'd3787208955;
	bram[953] <= 35'd3734821116;
	bram[954] <= 35'd3682425086;
	bram[955] <= 35'd3630012670;
	bram[956] <= 35'd3577600256;
	bram[957] <= 35'd3525171456;
	bram[958] <= 35'd3472742658;
	bram[959] <= 35'd3420297474;
	bram[960] <= 35'd3367852292;
	bram[961] <= 35'd3315390724;
	bram[962] <= 35'd3262929158;
	bram[963] <= 35'd3210451206;
	bram[964] <= 35'd3157973255;
	bram[965] <= 35'd3105487112;
	bram[966] <= 35'd3052992777;
	bram[967] <= 35'd3000490250;
	bram[968] <= 35'd2947979531;
	bram[969] <= 35'd2895460619;
	bram[970] <= 35'd2842941709;
	bram[971] <= 35'd2790406413;
	bram[972] <= 35'd2737871118;
	bram[973] <= 35'd2685327630;
	bram[974] <= 35'd2632784144;
	bram[975] <= 35'd2580224272;
	bram[976] <= 35'd2527664401;
	bram[977] <= 35'd2475096337;
	bram[978] <= 35'd2422528275;
	bram[979] <= 35'd2369943827;
	bram[980] <= 35'd2317359379;
	bram[981] <= 35'd2264774933;
	bram[982] <= 35'd2212174101;
	bram[983] <= 35'd2159573269;
	bram[984] <= 35'd2106972438;
	bram[985] <= 35'd2054363415;
	bram[986] <= 35'd2001746200;
	bram[987] <= 35'd1949120791;
	bram[988] <= 35'd1896503577;
	bram[989] <= 35'd1843869977;
	bram[990] <= 35'd1791236377;
	bram[991] <= 35'd1738602778;
	bram[992] <= 35'd1685960987;
	bram[993] <= 35'd1633311003;
	bram[994] <= 35'd1580661019;
	bram[995] <= 35'd1528011036;
	bram[996] <= 35'd1475352860;
	bram[997] <= 35'd1422694685;
	bram[998] <= 35'd1370028317;
	bram[999] <= 35'd1317361949;
	bram[1000] <= 35'd1264695582;
	bram[1001] <= 35'd1212021022;
	bram[1002] <= 35'd1159346463;
	bram[1003] <= 35'd1106663711;
	bram[1004] <= 35'd1053980959;
	bram[1005] <= 35'd1001298207;
	bram[1006] <= 35'd948615456;
	bram[1007] <= 35'd895924512;
	bram[1008] <= 35'd843233568;
	bram[1009] <= 35'd790542624;
	bram[1010] <= 35'd737851681;
	bram[1011] <= 35'd685152545;
	bram[1012] <= 35'd632453409;
	bram[1013] <= 35'd579754273;
	bram[1014] <= 35'd527055137;
	bram[1015] <= 35'd474356001;
	bram[1016] <= 35'd421656866;
	bram[1017] <= 35'd368949538;
	bram[1018] <= 35'd316242209;
	bram[1019] <= 35'd263543074;
	bram[1020] <= 35'd210835746;
	bram[1021] <= 35'd158128418;
	bram[1022] <= 35'd105421090;
	bram[1023] <= 35'd52713762;
end
endmodule
