/*
 * Copyright (C) 2014 Harmon Instruments, LLC
 *
 * This program is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with this program.  If not, see <http://www.gnu.org/licenses/
 *
 */

`timescale 1ns / 1ps

module sync_pulse(input ci, i, co, output reg o=0);
   reg it = 0;
   always @ (posedge ci)
     it <= i ^ it;
   wire it_o;
   sync sync_i(.c(co), .i(it), .o(it_o));
   reg 	it_o_prev = 0;
   always @ (posedge co)
     begin
	it_o_prev <= it_o;
	o <= it_o ^ it_o_prev;
     end
endmodule
/*
module sync_pulse_related(input ci, i, co, output reg o=0);
   reg it = 0;
   always @ (posedge ci)
     it <= it ^ i;
   reg 	it_prev = 0;
   always @ (posedge co)
     begin
	it_prev <= it;
	o <= it ^ it_prev;
     end
endmodule
*/
