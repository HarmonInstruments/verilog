module cosrom (
	input c, // clock
	input [9:0] a0, a1, // angle
	output [34:0] d0, d1);

wire [35:0] o0, o1;
assign d0 = o0[34:0];
assign d1 = o1[34:0];

RAMB36E1 #(
.DOA_REG(1),.DOB_REG(1),
.INIT_A(36'h000000000), .INIT_B(36'h000000000),
.RAM_MODE("TDP"),
.READ_WIDTH_A(36), .READ_WIDTH_B(36),
.WRITE_WIDTH_A(36), .WRITE_WIDTH_B(36),
.INIT_00(256'hFFE1A04AFFE9A040FFF08037FFF6002CFFFA6023FFFD6018FFFF400FFFFFE005),
.INIT_01(256'hFF752099FF87008FFF97A085FFA7007BFFB54072FFC24068FFCDE05DFFD86054),
.INIT_02(256'hFEB9A0E8FED560DEFEEFE0D4FF0920CAFF2140C1FF3800B6FF4DA0ADFF6200A3),
.INIT_03(256'hFDAF4137FDD4C12CFDF94124FE1C6119FE3E410FFE5F0106FE7E60FBFE9CA0F2),
.INIT_04(256'hFC55E185FC85617CFCB3A172FCE0A168FD0C615EFD370155FD60414AFD886141),
.INIT_05(256'hFAADE1D5FAE721CAFB1F41C1FB5621B7FB8BC1ADFBC021A3FBF34199FC254190),
.INIT_06(256'hF8B70223F8FA2219F93C2210F97CC205F9BC41FCF9FA81F2FA3781E8FA7341DE),
.INIT_07(256'hF6718272F6BE8268F70A425EF754C254F79E224BF7E62240F82D0237F872A22D),
.INIT_08(256'hF3DD62C0F43442B7F489C2ACF4DE22A3F5314299F583228FF5D3E286F623427B),
.INIT_09(256'hF0FAE30FF15B6304F1BAE2FCF21902F1F275E2E7F2D1A2DEF32C22D4F38562CA),
.INIT_0A(256'hEDC9E35DEE344353EE9D834AEF05633FEF6C2336EFD1A32CF035E322F0990319),
.INIT_0B(256'hEA4AA3ABEABEE3A2EB31C397EBA3838EEC140384EC83637BECF16370ED5E4367),
.INIT_0C(256'hE67D63FAE6FB43EFE77803E6E7F383DCE86DC3D2E8E6C3C8E95EA3BFE9D543B5),
.INIT_0D(256'hE2620447E2E9A43DE3702434E3F5642AE4796420E4FC4417E57DC40CE5FE2403),
.INIT_0E(256'hDDF8E495DE8A448BDF1A8482DFA96477E037246EE0C3C465E14F045AE1D92451),
.INIT_0F(256'hD94224E2D9DD44D9DA7724CFDB0FC4C5DBA744BCDC3D84B2DCD284A8DD66449E),
.INIT_10(256'hD43DE530D4E2A526D586451DD6288512D6C9A509D769A500D80864F6D8A5E4EC),
.INIT_11(256'hCEEC657DCF9AC573D048056AD0F40560D19EC556D248654DD2F0C543D397E539),
.INIT_12(256'hC94DE5CACA05E5C0CABCC5B7CB7265ADCC26C5A3CCDA059ACD8C0590CE3CC586),
.INIT_13(256'hC3628617C424260DC4E48603C5A3C5FAC661C5F0C71EA5E7C7DA45DDC894A5D3),
.INIT_14(256'hBD2A6663BDF5A65ABEBFA650BF886646C050063DC1166633C1DBA62AC29FA620),
.INIT_15(256'hB6A606AFB77AC6A6B84E469CB920A693B9F1C689BAC1C680BB908676BC5E066C),
.INIT_16(256'hAFD586FBB0B3C6F2B190C6E8B26CA6DFB34746D5B420C6CCB4F906C2B5D026B9),
.INIT_17(256'hA8B92747A9A0C73DAA874734AB6CA72BAC50C721AD33C718AE15870EAEF62705),
.INIT_18(256'hA1512793A2424789A332277FA420E776A50E876DA5FAE763A6E6275AA7D04751),
.INIT_19(256'h999DC7DD9A9867D59B91A7CA9C89E7C29D80E7B89E76A7AE9F6B67A6A05EC79B),
.INIT_1A(256'h919F882892A3681F93A6281694A7A80C95A8080396A747FA97A547F098A227E7),
.INIT_1B(256'h895688738A63C86A8B6FC8608C7AA8578D84684E8E8CE8448F94483B909A8832),
.INIT_1C(256'h80C328BD81D9A8B482EEE8AA840328A2851628988627E88E8738A8868848287C),
.INIT_1D(256'h77E5A907790568FE7A2408F57B4168EB7C5DA8E27D78C8D97E92A8CF7FAB88C7),
.INIT_1E(256'h6EBE89506FE78948710F493E7235E935735B492B747FA92375A2C91976C4C910),
.INIT_1F(256'h654E09996680299167B1098768E0C97E6A0F69756B3CE96C6C6949636D94895A),
.INIT_20(256'h5B9489E25CCFC9DA5E09C9D05F42A9C7607A69BE61B109B562E689AC641AE9A3),
.INIT_21(256'h51928A2B52D6AA215419CA19555BCA10569C8A0657DC49FE591AE9F55A5849EB),
.INIT_22(256'h47482A7348956A6A49E16A604B2C6A584C764A4F4DBF0A464F06AA3D504D2A34),
.INIT_23(256'h3CB5EABA3E0C2AB23F612AA840B52AA042080A974359AA8D44AA4A8545F9CA7C),
.INIT_24(256'h31DC6B02333B6AF834996AF035F64AE737520ADE38ACAAD53A064ACD3B5EAAC3),
.INIT_25(256'h26BBCB492823AB3F298A8B372AF04B2E2C54EB252DB86B1C2F1AEB14307C2B0A),
.INIT_26(256'h1B548B8E1CC54B861E34EB7D1FA38B752110EB6B227D4B6323E88B5A2552AB51),
.INIT_27(256'h0FA74BD51120CBCC12992BC314106BBA1586ABB216FBCBA9186FCBA019E2CB98),
.INIT_28(256'h03B42C1A05366C1206B78C0908378C0009B66BF70B344BEF0CB10BE60E2CABDD),
.INIT_29(256'hF77BEC5FF906CC57FA908C4EFC192C45FDA0AC3CFF272C3400ACAC2C0230EC22),
.INIT_2A(256'hEAFEECA3EC924C9BEE24AC93EFB5EC8AF1460C81F2D52C79F4632C70F5F00C67),
.INIT_2B(256'hDE3DACE7DFD98CDFE1746CD7E30E2CCEE4A6CCC5E63E6CBDE7D50CB5E96A8CAC),
.INIT_2C(256'hD138AD2BD2DCED22D4802D1AD6226D12D7C38D09D963AD01DB02CCF9DCA0CCF0),
.INIT_2D(256'hC3F04D6EC59CED65C748AD5EC8F34D55CA9CCD4CCC454D44CDECCD3CCF934D34),
.INIT_2E(256'hB6652DB1B81A2DA8B9CE2DA0BB812D98BD330D8FBEE3ED87C093CD7FC2428D76),
.INIT_2F(256'hA897CDF3AA550DEAAC114DE2ADCC8DDAAF86ADD1B13FEDCAB2F80DC1B4AF0DB8),
.INIT_30(256'h9A88AE349C4E2E2C9E128E239FD60E1CA1986E13A359CE0BA51A2E03A6D96DFA),
.INIT_31(256'h8C386E758E060E6D8FD28E64919E2E5D9368AE5495322E4C96FAAE4498C22E3C),
.INIT_32(256'h7DA78EB57F7D2EAD8151CEA583256E9D84F80E9586C9AE8D889A4E858A69CE7C),
.INIT_33(256'h6ED6AEF570B42EEC7290CEE5746C6EDD76470ED57820AECD79F94EC57BD0EEBD),
.INIT_34(256'h5FC62F3461ABAF2C63902F246573CF1D67564F146937CF0C6B186F056CF80EFD),
.INIT_35(256'h5076CF7252642F6B54508F63563BEF5B58264F535A0FCF4C5BF82F435DDFAF3C),
.INIT_36(256'h40E92FB042DE4FA944D26FA146C58F9948B7CF924AA8EF894C994F834E888F7A),
.INIT_37(256'h311DCFEE331A8FE635166FDF37114FD7390B2FCF3B040FC73CFC0FC03EF32FB9),
.INIT_38(256'h2115502B2319B023251D301C271F90132921300D2B21B0042D216FFE2F200FF5),
.INIT_39(256'h10D0506712DC305F14E7305816F1305018FA50491B0270411D09B03A1F0FF032),
.INIT_3A(256'h004F70A20262D09B047550940686D08C089750840AA6F07D0CB5B0760EC3706E),
.INIT_3B(256'hEF9370DDF1AE10D5F3C7F0CFF5E0D0C7F7F8D0C0FA0FD0B8FC25F0B1FE3B30AA),
.INIT_3C(256'hDE9CB117E0BEB110E2DFD109E5001102E71F50FAE93DB0F3EB5B30ECED77D0E5),
.INIT_3D(256'hCD6C3151CF955149D1BDB143D3E5113BD60BB135D831512DDA55F125DC79D11F),
.INIT_3E(256'hBC02518ABE329182C062117CC290B175C4BE516DC6EB1166C9171160CB421158),
.INIT_3F(256'hAA5FD1C2AC9731BBAECDB1B4B10351ADB33811A6B56BF19FB79EF198B9D11191),
.INIT_40(256'h988571F99AC3D1F39D0151EC9F3DD1E4A17991DEA3B471D7A5EE71D0A82791C9),
.INIT_41(256'h8673D23088B9122A8AFD72238D40F21C8F83921591C5520E9406320796465201),
.INIT_42(256'h742BB2667677B26078C2D2597B0D12527D56924C7F9F324581E6F23E842DD237),
.INIT_43(256'h61ADD29C640072956652528F68A352886AF372816D42D27B6F91527471DEF26D),
.INIT_44(256'h4EFAB2D15153F2CA53AC72C4560412BD585AD2B65AB0D2B05D05F2A95F5A52A3),
.INIT_45(256'h3C1333043E7312FF40D1F2F7433032F2458D72EA47EA12E54A45B2DD4CA092D7),
.INIT_46(256'h28F813372B5E53322DC3B32B30285325328C131E34EF13183751531239B2B30B),
.INIT_47(256'h15AA136A181693641A82535E1CED53581F57735121C0D34B242953442691333F),
.INIT_48(256'h0229D39C049C9396070E9390097FD38A0BF033830E5FD37D10CEB377133CD371),
.INIT_49(256'hEE7833CDF0F113C7F36933C1F5E093BBF85733B5FACCF3AEFD4213A9FFB653A2),
.INIT_4A(256'hDA95D3FDDD14D3F8DF92F3F1E21053EBE48D13E6E708F3DFE98413D9EBFE93D4),
.INIT_4B(256'hC683942DC9087427CB8C9421CE10141CD092B415D314940FD595B409D8163404),
.INIT_4C(256'hB242345BB4CCF456B756F450B9E0344ABC68D445BEF0943EC177B439C3FDF432),
.INIT_4D(256'h9DD2948AA062F483A2F2B47EA581D479A8101472AA9DB46DAD2A9467AFB6D462),
.INIT_4E(256'h893534B68BCB54B18E60D4AC90F574A5938994A1961CD49A98AF74959B41548F),
.INIT_4F(256'h746B34E37706D4DD79A1D4D87C3C34D37ED5B4CC816EB4C88406D4C1869E74BD),
.INIT_50(256'h5F75350F6216550964B6B503675694FF69F594F86C9414F46F31B4ED71CED4E9),
.INIT_51(256'h4A53F5394CFA75344FA0552F5245752954E9F524578DB51E5A30D5195CD35514),
.INIT_52(256'h3508756337B4355E3A5F55593D09B5533FB3754E425C95494505154447ACD53E),
.INIT_53(256'h1F93758C2244558724F4958227A4157C2A5315782D0175732FAF156D325C1568),
.INIT_54(256'h09F5B5B40CAB95AF0F60D5AA121595A614C995A0177CF59B1A2FD5971CE1F591),
.INIT_55(256'hF43015DCF6EAF5D7F9A535D2FC5ED5CDFF17D5C801D035C30487F5BE073F35BA),
.INIT_56(256'hDE437602E10335FEE3C235F8E680B5F4E93E95EFEBFBD5EAEEB895E6F17495E0),
.INIT_57(256'hC830B628CAF51623CDB8F61FD07C1619D33ED616D600D610D8C2560CDB833607),
.INIT_58(256'hB1F8964DB4C19648B78A1644BA51F63FBD19363ABFDFF636C2A61631C56BB62D),
.INIT_59(256'h9B9BF6719E69766CA1367668A402D663A6CEB65FA99A165BAC64D656AF2EF651),
.INIT_5A(256'h851BB69487EDB6908ABF168B8D8FF68790603682932FF67E95FF367A98CDD675),
.INIT_5B(256'h6E78D6B6714F16B27424B6AD76F9F6AA79CE96A57CA2B6A17F76369C82493698),
.INIT_5C(256'h57B3F6D75A8E76D45D6856CF6041B6CB631A96C765F2F6C368CAB6BE6BA216BB),
.INIT_5D(256'h40CE36F843ACB6F4468AB6F0496836EC4C4536E84F2196E351FD96E054D916DC),
.INIT_5E(256'h29C857182CAAB7132F8CB710326E370C354F3708382FB7043B0FB7003DEF36FC),
.INIT_5F(256'h12A3373715897732186F572F1B54B72B1E399727211DF7232401D71F26E5571C),
.INIT_60(256'hFB5FB754FE49B7500133574D041C77490705374609ED57410CD5173E0FBC573A),
.INIT_61(256'hE3FED771E6EC776DE9D9B76AECC69767EFB2D762F29ED760F58A375BF8753758),
.INIT_62(256'hCC81778DCF729789D2635786D553B783D843977FDB33177CDE221778E110B775),
.INIT_63(256'hB4E857A8B7DCF7A5BAD137A2BDC4F79EC0B8579BC3AB3797C69DB794C98FD791),
.INIT_64(256'h9D3497C2A02C97C0A323F7BBA61B17B9A911D7B6AC0817B2AEFDF7AFB1F357AB),
.INIT_65(256'h856717DC886237D98B5CD7D58E5717D29150F7CF944A77CC974397C99A3C57C6),
.INIT_66(256'h6D80B7F5707ED7F1737C97EE7679F7EB7976F7E87C7397E57F6FB7E1826B97DF),
.INIT_67(256'h5582380B588358095B8418065E847803618457FF6483F7FD678337FA6A8217F7),
.INIT_68(256'h3D6CD8224070B81F4374581D46777819497A58174C7CD8144F7F18125280D80E),
.INIT_69(256'h254158382847F8352B4E38322E5438303159B82C345F182B3763F8273A689825),
.INIT_6A(256'h0D00984C1009D84A1312B847161B5845192398421C2B783F1F33183D223A583A),
.INIT_6B(256'hF4AB9860F7B7585EFAC2B85BFDCDD85900D8985603E3185406ED385109F7184F),
.INIT_6C(256'hDC435872DF517871E25F386EE56CB86CE879D869EB86B867EE935865F19F9862),
.INIT_6D(256'hC3C8D885C6D91882C9E91880CCF8D87ED008587CD3177879D6267878D9351875),
.INIT_6E(256'hAB3CB895AE4F3894B1615891B473388FB784D88DBA96388BBDA75889C0B83887),
.INIT_6F(256'h92A038A595B4B8A498C8D8A19BDCD8A09EF0789DA203F89CA5171899A82A1898),
.INIT_70(256'h79F438B47D0A98B3802098B0833678AF864C18AD896178AB8C76B8AA8F8B98A7),
.INIT_71(256'h613998C26451B8C1676998BF6A8138BD6D98B8BC70AFF8BA73C6F8B876DDB8B6),
.INIT_72(256'h487178D04B8B38CE4EA4B8CC51BE18CB54D738C957F018C75B08D8C65E2158C4),
.INIT_73(256'h2F9C98DC32B7D8DA35D2F8D938EDD8D73C0878D53F2318D5423D58D2455778D1),
.INIT_74(256'h16BBF8E719D898E51CF538E5201178E2232DB8E22649B8E0296578DE2C8118DD),
.INIT_75(256'hFDD098F100EE98F0040C78EF072A18ED0A4798EC0D64F8EB108218E9139F18E8),
.INIT_76(256'hE4DB98FBE7FAB8F9EB19B8F8EE3898F7F15738F5F475D8F5F79438F3FAB278F2),
.INIT_77(256'hCBDD9902CEFDD902D21DD900D53DD900D85D98FEDB7D58FEDE9CD8FCE1BC38FB),
.INIT_78(256'hB2D7D90AB5F8F909B919F908BC3AD907BF5B9906C27C5906C59CD904C8BD5904),
.INIT_79(256'h99CB19109CED1910A00ED90EA330990EA652390DA973D90DAC95390BAFB6990B),
.INIT_7A(256'h80B8791583DB191586FDB9158A2019138D4279139064D9139386F91196A91911),
.INIT_7B(256'h67A0F91A6AC419196DE73919710A5919742D3917775039187A7319177D95D916),
.INIT_7C(256'h4E85591D51A8F91D54CC991D57F0191C5B13991C5E36F91B615A591B647DB91B),
.INIT_7D(256'h3566B920388AB9203BAE991F3ED2791F41F6591F451A391F483DF91E4B61B91E),
.INIT_7E(256'h1C4619211F6A3921228E592125B2792128D699212BFAB9212F1EB9203242B920),
.INIT_7F(256'h0324592206489922096CD9220C9119220FB5592212D9792115FDB9221921F922),
.INITP_00(256'h7777777777777777777777777777777777777777777777777777777777777777),
.INITP_01(256'h7777777777777777777777777777777777777777777777777777777777777777),
.INITP_02(256'h7777777777777777777777777777777777777777777777777777777777777777),
.INITP_03(256'h7777777777777777777777777777777777777777777777777777777777777777),
.INITP_04(256'h7777777777777777777777777777777777777777777777777777777777777777),
.INITP_05(256'h6666666666666666666666666666666666666666666666666666667777777777),
.INITP_06(256'h6666666666666666666666666666666666666666666666666666666666666666),
.INITP_07(256'h5555555555555555555555555555555555555555666666666666666666666666),
.INITP_08(256'h5555555555555555555555555555555555555555555555555555555555555555),
.INITP_09(256'h4444444444444444444444444444444444444444444444444444444455555555),
.INITP_0A(256'h3333333333333333333334444444444444444444444444444444444444444444),
.INITP_0B(256'h3333333333333333333333333333333333333333333333333333333333333333),
.INITP_0C(256'h2222222222222222222222222222222222222222222222222222222222333333),
.INITP_0D(256'h1111111111111111111111111111111111112222222222222222222222222222),
.INITP_0E(256'h0000000000000000011111111111111111111111111111111111111111111111),
.INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
.SIM_DEVICE("7SERIES"))
RAMB36E1_inst (
.CASCADEOUTA(), .CASCADEOUTB(),
.DBITERR(), .ECCPARITY(), .RDADDRECC(), .SBITERR(),
.DOADO(o0[31:0]),
.DOPADOP(o0[35:32]),
.DOBDO(o1[31:0]),
.DOPBDOP(o1[35:32]),
.CASCADEINA(1'b0), .CASCADEINB(1'b0),
.INJECTDBITERR(1'b0), .INJECTSBITERR(1'b0),
.ADDRARDADDR({1'b0,a0,5'd0}),
.CLKARDCLK(c),
.ENARDEN(1'b1),
.REGCEAREGCE(1'b1),
.RSTRAMARSTRAM(1'b0),
.RSTREGARSTREG(1'b0),
.WEA(4'b0),
.DIADI(32'h0),
.DIPADIP(4'h0),
.ADDRBWRADDR({1'b0,a1,5'd0}),
.CLKBWRCLK(c),
.ENBWREN(1'b1),
.REGCEB(1'b1),
.RSTRAMB(1'b0),
.RSTREGB(1'b0),
.WEBWE(8'b0),
.DIBDI(32'h0),
.DIPBDIP(4'h0));
endmodule
